//module DrawPlayer(
//	input [4:0] x , 
//	input [3:0] y ,
//	input [1:0] behavior,
//	input direction ,
//	input [1:0] period ,
//	input Draw_En,
//
//
//)
//
//
//
//
//
//endmodule
