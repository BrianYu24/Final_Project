//module DrawEnemy(
//	input [4:0] x [5], 
//	input [3:0] y [5],
//	input [2:0] Count,
//	input [1:0] behavior [5],
//	input direction [5],
//	input [1:0] period [5],
//	input Draw_En,
//
//
//)
//
//
//
//
//
//endmodule
